/*
 * Module: register_file
 *
 * Description: Branch control logic. Only sets the branch control bits based on the
 * branch instruction
 *
 * Inputs:
 * 1) clk
 * 2) reset signal rst
 * 3) 5-bit rs1 address rs1_i
 * 4) 5-bit rs2 address rs2_i
 * 5) 5-bit rd address rd_i
 * 6) DWIDTH-wide data writeback datawb_i
 * 7) register write enable regwren_i
 * Outputs:
 * 1) 32-bit rs1 data rs1data_o
 * 2) 32-bit rs2 data rs2data_o
 */

module register_file(
  input  logic        clk_i,
  input  logic        reset_i,
  input  logic [4:0]  rs1_i,
  input  logic [4:0]  rs2_i,
  input  logic [4:0]  rd_i,
  input  logic        regwren_i,
  input  logic [31:0] datawb_i,
  output logic [31:0] rs1_data_o,
  output logic [31:0] rs2_data_o
);
  logic [31:0] regs [31:0];
  integer i;

  // Combinational reads
  assign rs1_data_o = (rs1_i == 5'd0) ? 32'd0 : regs[rs1_i];
  assign rs2_data_o = (rs2_i == 5'd0) ? 32'd0 : regs[rs2_i];

  always_ff @(posedge clk_i) begin
    if (reset_i) begin
      for (i = 0; i < 32; i++) regs[i] <= 32'd0;
      regs[5'd2] <= 32'h4000_0002;  // Seed x2
    end else if (regwren_i && (rd_i != 5'd0)) begin
      regs[rd_i] <= datawb_i;
    end
  end
endmodule
