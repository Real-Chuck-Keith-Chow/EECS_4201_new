// ----  Probes  ----
`define PROBE_ADDR      f_pc      //connection where pc_o and addr_i meet
`define PROBE_DATA_IN   data_i    //input for data in memory
`define PROBE_DATA_OUT  data_o    //output for data in memory
`define PROBE_READ_EN   read_en   
`define PROBE_WRITE_EN  write_en  

`define PROBE_F_PC      f_pc    //input memory address/PC 
`define PROBE_F_INSN    f_inst  //fetch_insn_o 

// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----

