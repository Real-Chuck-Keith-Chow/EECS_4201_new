/*
 * Good practice to define constants and refer to them in the
 * design files. An example of some constants are provided to you
 * as a starting point
 *
 */
`ifndef CONSTANTS_SVH_
`define CONSTANTS_SVH_

parameter logic [31:0] ZERO = 32'd0;
parameter logic [31:0] SP_RESET = 32'h0110_0000;

/*
 * Define constants as required...
 */

`endif
