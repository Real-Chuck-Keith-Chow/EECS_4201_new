/*
 * Module: pd2
 *
 * Description: Top level module that will contain sub-module instantiations.
 *
 * Inputs:
 * 1) clk
 * 2) reset signal
 */

module pd2 #(
    parameter int AWIDTH = 32,
    parameter int DWIDTH = 32)(
    input logic clk,
    input logic reset
);


    control #()control1();
    decode #()decode1();
    igen #()igen1();
    memory #()memory1();
    
    
 /*
  * Instantiate other submodules and
  * probes. To be filled by student...
  *
  */

endmodule : pd2
