
`define PROBE_F_PC           PROBE_F_PC_q
`define PROBE_F_INSN         PROBE_F_INSN_q

`define PROBE_D_PC           PROBE_D_PC_q
`define PROBE_D_OPCODE       D_opcode
`define PROBE_D_RD           D_rd
`define PROBE_D_FUNCT3       D_funct3
`define PROBE_D_RS1          D_rs1
`define PROBE_D_RS2          D_rs2
`define PROBE_D_FUNCT7       D_funct7
`define PROBE_D_IMM          PROBE_D_IMM_q
`define PROBE_D_SHAMT        D_shamt

`define PROBE_R_WRITE_ENABLE      PROBE_R_WE_q
`define PROBE_R_WRITE_DESTINATION PROBE_R_RD_q
`define PROBE_R_WRITE_DATA        PROBE_R_WD_q
`define PROBE_R_READ_RS1          PROBE_R_RS1_q
`define PROBE_R_READ_RS2          PROBE_R_RS2_q
`define PROBE_R_READ_RS1_DATA     PROBE_R_RS1D_q
`define PROBE_R_READ_RS2_DATA     PROBE_R_RS2D_q

`define PROBE_E_PC                PROBE_E_PC_q
`define PROBE_E_ALU_RES           PROBE_E_ALU_q
`define PROBE_E_BR_TAKEN          PROBE_E_TAKEN_q

`define PROBE_M_PC                PROBE_M_PC_q
`define PROBE_M_ADDRESS           PROBE_M_ADDR_q
`define PROBE_M_SIZE_ENCODED      PROBE_M_SIZE_q
`define PROBE_M_DATA              PROBE_M_DATA_q

`define PROBE_W_PC                PROBE_W_PC_q
`define PROBE_W_ENABLE            PROBE_W_EN_q
`define PROBE_W_DESTINATION       PROBE_W_DEST_q
`define PROBE_W_DATA              PROBE_W_DATA_q

// ----  Top module  ----
`define TOP_MODULE  pd4
// ----  Top module  ----
