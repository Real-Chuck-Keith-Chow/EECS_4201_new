`include "constants.svh"
